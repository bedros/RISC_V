`define BYTE 2'b00
`define WORD 2'b01
`define DWORD 2'b10

//不支持非对齐字节读写
//非对齐读写将会产生异常

module BIU(
);
endmodule
